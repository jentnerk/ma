/usr/pack/gf-45soi-kgf/dz/../gf/45RFSOI-RF/V1.0_1.1/PlaceRoute/Innovus/lef/45RFSOI_8LM_3Mx_1Cx_1Ux_2Ox_LD_tech.lef