/usr/pack/gf-45soi-kgf/arm/gf/45rfsoi/sc9_base_uvt/r0p0/lef/sc9_soi12s0_base_uvt.lef