/usr/pack/gf-45soi-kgf/arm/gf/45rfsoi/sc9_base_hvt/r0p0/lef/sc9_soi12s0_base_hvt.lef